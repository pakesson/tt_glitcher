`default_nettype none

module uart_handler #(
    parameter CLK_FREQ = 50_000_000,
    parameter BAUD_RATE = 115200
) (
    input wire        rst,
    input wire        clk,
    input wire        uart_rx_i,
    output wire       uart_tx_o,
    output reg [15:0] delay_o,
    output reg [7:0]  width_o,
    output reg [7:0]  num_pulses_o,
    output reg [15:0] pulse_spacing_o,
    output reg        pulse_en_o,
    output reg        reset_en_o,
    output reg [15:0] reset_length_o
);

    wire uart_rx_valid;
    wire [7:0] uart_rx_data;
    
    uart_rx #(
        .CLK_FREQ(CLK_FREQ),
        .BAUD_RATE(BAUD_RATE)
    ) rxi (
        .clk(clk),
        .rst(rst),
        .rx_i(uart_rx_i),
        .data_o(uart_rx_data),
        .data_valid_o(uart_rx_valid)
    );

    wire uart_tx_busy;
    wire uart_tx_rdy = !uart_tx_busy;
    reg uart_tx_en;
    reg [7:0] uart_tx_data;

    uart_tx #(
        .CLK_FREQ(CLK_FREQ),
        .BAUD_RATE(BAUD_RATE)
    ) txi (
        .clk(clk),
        .rst(rst),
        .tx_data_i(uart_tx_data),
        .tx_enable_i(uart_tx_en),
        .tx_o(uart_tx_o),
        .tx_busy_o(uart_tx_busy)
    );

    reg [3:0] state;
    localparam STATE_IDLE = 4'd0;
    localparam STATE_DELAY1 = 4'd2;
    localparam STATE_DELAY0 = 4'd3;
    localparam STATE_WIDTH = 4'd4;
    localparam STATE_NUM_PULSES = 4'd5;
    localparam STATE_PULSE_SPACING1 = 4'd6;
    localparam STATE_PULSE_SPACING0 = 4'd7;
    localparam STATE_RESET_LENGTH1 = 4'd8;
    localparam STATE_RESET_LENGTH0 = 4'd9;
    localparam STATE_TRIGGER_PULSE = 4'd10;
    localparam STATE_SEND_HELLO = 4'd11;

    reg [2:0] hello_state;

    always @(posedge clk) begin
        if (rst) begin
            delay_o <= 16'd0;
            width_o <= 8'd0;
            num_pulses_o <= 8'd0;
            pulse_spacing_o <= 16'd0;
            pulse_en_o <= 1'b0;
            reset_en_o <= 1'b0;
            reset_length_o <= 16'd0;

            uart_tx_en <= 1'b0;
            uart_tx_data <= 8'd0;

            state <= STATE_IDLE;
            hello_state <= 3'd0;
        end else begin
            uart_tx_en <= 1'b0;
            pulse_en_o <= 1'b0;
            reset_en_o <= 1'b0;

            case(state)
                STATE_IDLE:
                    if (uart_rx_valid) begin
                        case (uart_rx_data)
                            8'h64: state <= STATE_DELAY1;         // 'd'
                            8'h77: state <= STATE_WIDTH;          // 'w'
                            8'h6E: state <= STATE_NUM_PULSES;     // 'n'
                            8'h73: state <= STATE_PULSE_SPACING1; // 's'
                            8'h72: state <= STATE_RESET_LENGTH1;  // 'r'
                            8'h74: state <= STATE_TRIGGER_PULSE;  // 't'
                            8'h68: state <= STATE_SEND_HELLO;     // 'h'
                            default: 
                                state <= STATE_IDLE;
                        endcase
                    end
                STATE_DELAY1:
                    if (uart_rx_valid) begin
                        delay_o[15:8] <= uart_rx_data;
                        state <= STATE_DELAY0;
                    end
                STATE_DELAY0:
                    if (uart_rx_valid) begin
                        delay_o[7:0] <= uart_rx_data;
                        state <= STATE_IDLE;
                    end
                STATE_WIDTH:
                    if (uart_rx_valid) begin
                        width_o <= uart_rx_data;
                        state <= STATE_IDLE;
                    end
                STATE_NUM_PULSES:
                    if (uart_rx_valid) begin
                        num_pulses_o <= uart_rx_data;
                        state <= STATE_IDLE;
                    end
                STATE_PULSE_SPACING1:
                    if (uart_rx_valid) begin
                        pulse_spacing_o[15:8] <= uart_rx_data;
                        state <= STATE_PULSE_SPACING0;
                    end
                STATE_PULSE_SPACING0:
                    if (uart_rx_valid) begin
                        pulse_spacing_o[7:0] <= uart_rx_data;
                        state <= STATE_IDLE;
                    end
                STATE_RESET_LENGTH1:
                    if (uart_rx_valid) begin
                        reset_length_o[15:8] <= uart_rx_data;
                        state <= STATE_RESET_LENGTH0;
                    end
                STATE_RESET_LENGTH0:
                    if (uart_rx_valid) begin
                        reset_length_o[7:0] <= uart_rx_data;
                        state <= STATE_IDLE;
                    end
                STATE_TRIGGER_PULSE:
                    begin
                        if (reset_length_o != 16'd0)
                            // Set reset_en high for one clock cycle
                            reset_en_o <= 1'b1;
                        else
                            // Set pulse_en high for one clock cycle
                            pulse_en_o <= 1'b1;
                        state <= STATE_IDLE;
                    end
                STATE_SEND_HELLO:
                    if (uart_tx_rdy && !uart_tx_en) begin
                        case (hello_state)
                            3'd0: begin
                                uart_tx_data <= 8'h48;
                                uart_tx_en <= 1'b1;
                                hello_state <= 3'd1;
                            end
                            3'd1: begin
                                uart_tx_data <= 8'h65;
                                uart_tx_en <= 1'b1;
                                hello_state <= 3'd2;
                            end
                            3'd2: begin
                                uart_tx_data <= 8'h6C;
                                uart_tx_en <= 1'b1;
                                hello_state <= 3'd3;
                            end
                            3'd3: begin
                                uart_tx_data <= 8'h6C;
                                uart_tx_en <= 1'b1;
                                hello_state <= 3'd4;
                            end
                            3'd4: begin
                                uart_tx_data <= 8'h6F;
                                uart_tx_en <= 1'b1;
                                hello_state <= 3'd5;
                            end
                            3'd5: begin
                                uart_tx_data <= 8'h0A;
                                uart_tx_en <= 1'b1;
                                hello_state <= 3'd0;
                                state <= STATE_IDLE;
                            end
                            default:
                                begin
                                    hello_state <= 3'd0;
                                    state <= STATE_IDLE;
                                end
                        endcase
                    end
                default:
                    state <= STATE_IDLE;
            endcase
        end
    end

endmodule